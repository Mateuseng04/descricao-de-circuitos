library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity subtrator4bits is
    port (
        a, b      : in  std_logic_vector(3 downto 0);
        resultado : out std_logic_vector(3 downto 0);
        borrow    : out std_logic
    );
end subtrator4bits;

architecture comportamento of subtrator4bits is

    signal a_ext, b_ext : signed(4 downto 0);
    signal sub_tmp      : signed(4 downto 0);

begin

    a_ext <= signed('0' & a);  
    b_ext <= signed('0' & b);

    sub_tmp <= a_ext - b_ext;

    resultado <= std_logic_vector(sub_tmp(3 downto 0));

    borrow <= '1' when unsigned(a) < unsigned(b) else '0';

end comportamento;
